`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
//////////////////////////////////////////////////////////////////////////////////


package common;
typedef enum {
    S0,
    S1,
    S2,
    S3,
    S4
} example_states;

endpackage
